# 
# +++++++++++++++++++++++++++++++++++++++++++++
# ++++++++++     DESIGN HIERARCHY    ++++++++++
# +++++++++++++++++++++++++++++++++++++++++++++
# 
# 
# CUMULATIVE SUMMARY
# =============================================
# |    Coverage Type    | Weight | Hits/Total |
# =============================================
# | Covergroup Coverage |      1 |    56.250% |
# |---------------------|--------|------------|
# | Types               |        |      0 / 1 |
# =============================================
# CUMULATIVE INSTANCE-BASED COVERAGE: 56.250%
# COVERED INSTANCES: 0 / 1
# FILES: 1
# 
# 
# INSTANCE - /tb : work.tb
# 
# 
#     SUMMARY
#     ==========================================================================
#     |    Coverage Type    | Weight | Local Hits/Total | Recursive Hits/Total |
#     ==========================================================================
#     | Covergroup Coverage |      1 |          56.250% |              56.250% |
#     |---------------------|--------|------------------|----------------------|
#     | Types               |        |            0 / 1 |                0 / 1 |
#     ==========================================================================
#     WEIGHTED AVERAGE LOCAL: 56.250%
#     WEIGHTED AVERAGE RECURSIVE: 56.250%
# 
# 
#     COVERGROUP COVERAGE
#     =================================================
#     |  Covergroup  |  Hits   |  Goal /  |  Status   |
#     |              |         | At Least |           |
#     =================================================
#     | TYPE /tb/c_g | 56.250% | 100.000% | Uncovered |
#     =================================================
# 
# 
# +++++++++++++++++++++++++++++++++++++++++++++
# ++++++++++       DESIGN UNITS      ++++++++++
# +++++++++++++++++++++++++++++++++++++++++++++
# 
# 
# CUMULATIVE SUMMARY
# =============================================
# |    Coverage Type    | Weight | Hits/Total |
# =============================================
# | Covergroup Coverage |      1 |    56.250% |
# |---------------------|--------|------------|
# | Types               |        |      0 / 1 |
# =============================================
# CUMULATIVE DESIGN-BASED COVERAGE: 56.250%
# COVERED DESIGN UNITS: 0 / 1
# FILES: 1
# 
# 
# MODULE - work.tb
# 
# 
#     SUMMARY
#     =============================================
#     |    Coverage Type    | Weight | Hits/Total |
#     =============================================
#     | Covergroup Coverage |      1 |    56.250% |
#     |---------------------|--------|------------|
#     | Types               |        |      0 / 1 |
#     =============================================
#     WEIGHTED AVERAGE: 56.250%
# 
# 
#     COVERGROUP COVERAGE
#     =================================================
#     |  Covergroup  |  Hits   |  Goal /  |  Status   |
#     |              |         | At Least |           |
#     =================================================
#     | TYPE /tb/c_g | 56.250% | 100.000% | Uncovered |
#     =================================================
# 
exit
# VSIM: Simulation has finished.
Done
