Uploading......!
